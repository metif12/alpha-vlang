module main

fn main() {
	println('Starting...')

	log := parse() ?

	println(log)
}
