module main

[heap]
struct Place {
	inputs []string
	outputs []string
}