module main

import time

[heap]
struct Event {
	id        string
	title     string
	timestamp time.Time
}
